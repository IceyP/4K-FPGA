module s7_box(                                                         
	A                           ,                                      
	SPO                                                               
	);                                                                 
                                                                       
input   [5:0]                   A                                   ;  
output  [3:0]                   SPO                                 ;  

assign  SPO = (A==6'h00) ? 4'b0100:
              (A==6'h01) ? 4'b1101:
              (A==6'h02) ? 4'b1011:
              (A==6'h03) ? 4'b0000:
              (A==6'h04) ? 4'b0010:
              (A==6'h05) ? 4'b1011:
              (A==6'h06) ? 4'b1110:
              (A==6'h07) ? 4'b0111:
              (A==6'h08) ? 4'b1111:
              (A==6'h09) ? 4'b0100:
              (A==6'h0A) ? 4'b0000:
              (A==6'h0B) ? 4'b1001:
              (A==6'h0C) ? 4'b1000:
              (A==6'h0D) ? 4'b0001:
              (A==6'h0E) ? 4'b1101:
              (A==6'h0F) ? 4'b1010:
              (A==6'h10) ? 4'b0011:
              (A==6'h11) ? 4'b1110:
              (A==6'h12) ? 4'b1100:
              (A==6'h13) ? 4'b0011:
              (A==6'h14) ? 4'b1001:
              (A==6'h15) ? 4'b0101:
              (A==6'h16) ? 4'b0111:
              (A==6'h17) ? 4'b1100:
              (A==6'h18) ? 4'b0101:
              (A==6'h19) ? 4'b0010:
              (A==6'h1A) ? 4'b1010:
              (A==6'h1B) ? 4'b1111:
              (A==6'h1C) ? 4'b0110:
              (A==6'h1D) ? 4'b1000:
              (A==6'h1E) ? 4'b0001:
              (A==6'h1F) ? 4'b0110:
              (A==6'h20) ? 4'b0001:
              (A==6'h21) ? 4'b0110:
              (A==6'h22) ? 4'b0100:
              (A==6'h23) ? 4'b1011:
              (A==6'h24) ? 4'b1011:
              (A==6'h25) ? 4'b1101:
              (A==6'h26) ? 4'b1101:
              (A==6'h27) ? 4'b1000:
              (A==6'h28) ? 4'b1100:
              (A==6'h29) ? 4'b0001:
              (A==6'h2A) ? 4'b0011:
              (A==6'h2B) ? 4'b0100:
              (A==6'h2C) ? 4'b0111:
              (A==6'h2D) ? 4'b1010:
              (A==6'h2E) ? 4'b1110:
              (A==6'h2F) ? 4'b0111:
              (A==6'h30) ? 4'b1010:
              (A==6'h31) ? 4'b1001:
              (A==6'h32) ? 4'b1111:
              (A==6'h33) ? 4'b0101:
              (A==6'h34) ? 4'b0110:
              (A==6'h35) ? 4'b0000:
              (A==6'h36) ? 4'b1000:
              (A==6'h37) ? 4'b1111:
              (A==6'h38) ? 4'b0000:
              (A==6'h39) ? 4'b1110:
              (A==6'h3A) ? 4'b0101:
              (A==6'h3B) ? 4'b0010:
              (A==6'h3C) ? 4'b1001:
              (A==6'h3D) ? 4'b0011:
              (A==6'h3E) ? 4'b0010:
              (A==6'h3F) ? 4'b1100:
			  4'b1100;
endmodule